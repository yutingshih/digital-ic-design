module Token;

parameter ZERO = 5'h0;
parameter ONE = 5'h1;
parameter TWO = 5'h2;
parameter THREE = 5'h3;
parameter FOUR = 5'h4;
parameter FIVE = 5'h5;
parameter SIX = 5'h6;
parameter SEVEN = 5'h7;
parameter EIGHT = 5'h8;
parameter NINE = 5'h9;
parameter TEN = 5'ha;
parameter ELEVEN = 5'hb;
parameter TWELVE = 5'hc;
parameter THIRTEEN = 5'hd;
parameter FOURTEEN = 5'he;
parameter FIFTEEN = 5'hf;

parameter LEFT  = 5'h18;  // (
parameter RIGHT = 5'h19;  // )
parameter MUL   = 5'h1a;  // *
parameter ADD   = 5'h1b;  // +
parameter SUB   = 5'h1d;  // -
parameter EVAL  = 5'h1f;  // =

parameter UNKNOWN = 'bx;

endmodule
