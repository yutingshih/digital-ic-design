module Constants;

parameter BIAS = 13'h1FF4;
parameter KERN0 = 13'h1FFF;
parameter KERN1 = 13'h1FFE;
parameter KERN2 = 13'h1FFF;
parameter KERN3 = 13'h1FFC;
parameter KERN4 = 13'h0010;
parameter KERN5 = 13'h1FFC;
parameter KERN6 = 13'h1FFF;
parameter KERN7 = 13'h1FFE;
parameter KERN8 = 13'h1FFF;

endmodule
